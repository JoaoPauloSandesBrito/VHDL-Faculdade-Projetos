library verilog;
use verilog.vl_types.all;
entity ula4b_vlg_vec_tst is
end ula4b_vlg_vec_tst;
